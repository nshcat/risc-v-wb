`ifndef _WB_BUS_H
`define _WB_BUS_H

`endif