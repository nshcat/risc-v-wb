module top(
    input logic clk_in,
    input logic rst_in
);

endmodule
