`ifndef _CORE_DEFINES_H
`define _CORE_DEFINES_H



`endif